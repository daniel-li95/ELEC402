/ubc/ece/home/ugrads/v/v6d9/ELEC402/Modelsim_50995133/ELEC402/PnR/in/gsclib045_macro.lef